//
//
//
//`define NUM_SPRITE_REGS 10
////module player_mapper (  input [24:0] sprite_info,
////                        input Clk,
////                        input [9:0] DrawX, DrawY,
////                        output logic [3:0] palette_out);
////
////
////    /*-- Mapping from the sprite list to variables--*/
////    //logic [4:0] sprite_idx;
////    logic [8:0] XCoord;
////    logic [9:0] YCoord;
////    logic sprite_en, draw_sprite;
////    assign XCoord = sprite_info[18:10];
////    assign YCoord = sprite_info[9:0];
////    assign sprite_en = sprite_info[19];
////    
////    
////    /*-- Calculate all boundaries, x/y coord is top left --*/
////    int leftBound, rightBound, topBound, lowerBound;
////    
////    assign leftBound = XCoord;
////    assign rightBound = XCoord+31;
////    assign topBound = YCoord;
////    assign lowerBound = YCoord+47;
////
////    /*-- Check if DrawX/DrawY is within boundaries, check if I should draw the sprite --*/
////    always_comb begin
////        if (DrawX>=leftBound & DrawX<=rightBound & sprite_en
////            & DrawY>=lowerBound & DrawY<=topBound) begin
////                draw_sprite = 1'b1;
////            end else begin
////                draw_sprite = 1'b0;
////            end
////    end
////
////    /*-- Calculate the pixel access index (to access the rom) --*/
////    int Xsprite, Ysprite, xOffset, yOffset, pixel_access;
////    assign Xsprite = leftBound - XCoord;
////    assign Ysprite = topBound - YCoord;
////    assign xOffset = Xsprite >> 5;
////    assign pixel_access = (32*Ysprite)+xOffset;
////
////    logic [3:0] palette_idx, data_in;
////
////    playerCenterROM player(.data_in(4'b0), .write_address(11'b0), .read_address(pixel_access), .we(1'b0), .Clk(Clk), .data_out(palette_idx));
////    
////    assign palette_out = (draw_sprite) ? palette_idx : 4'b0;
////    
////
////endmodule
//
//
//// this module takes drawX, drawY coordinates and outputs the RGB data to be used
//module color_mapper (   input Clk, Reset,
//                        input [9:0] DrawX, DrawY,
//                        output logic [3:0] palette_out );
//
//    
//    /*-- Registers hold the encoding for each sprite --*/
//    // X/Y coordinates should be edited in software
//    // encoding: [24:20] sprite_idx, [19] enable, [18:10] xcoord, [9:0] y coord
//    // order: player_center[0], winged_eye[1], enemy_ghost[2], enemy_fairy[3], bullet[4] 
//
//    /*-- color data for each sprite. Need to process to choose which to use --*/
//    logic [3:0] playerColor, wEyeColor, ghostColor, fairyColor, bulletColor, outputColor;
//
//    /*-- These modules provide color data based on whether each individual sprite should be printed --*/
//    player_mapper player1 (.sprite_info(20'h88020), .Clk(Clk), .DrawX(DrawX), .DrawY(DrawY), .palette_out(playerColor));
////	 player_mapper player1 (.sprite_info(SPRITE_REGS[0]), .Clk(Clk), .DrawX(DrawX), .DrawY(DrawY), .palette_out(playerColor));
////    winged_eye eye1 (.sprite_info(SPRITE_REGS[1]), .Clk(Clk), .DrawX(DrawX), .DrawY(DrawY), .palette_out(wEyeColor));
////    enemy_ghost ghost1 (.sprite_info(SPRITE_REGS[2]), .Clk(Clk), .DrawX(DrawX), .DrawY(DrawY), .palette_out(ghostColor));
////    enemy_fairy fairy1 (.sprite_info(SPRITE_REGS[3]), .Clk(Clk), .DrawX(DrawX), .DrawY(DrawY), .palette_out(fairyColor));
////    bullet b1 (.sprite_info(SPRITE_REGS[4]), .Clk(Clk), .DrawX(DrawX), .DrawY(DrawY), .palette_out(bulletColor));
//
//    /*-- Process the color data from each sprite, if statements in priority to be set --*/
//    always_comb begin
////        if (playerColor!=0)
////            outputColor = playerColor;
////        else if (wEyeColor!=0)
////            outputColor = wEyeColor;
////        else if (ghostColor!=0)
////            outputColor = ghostColor;
////        else if (fairyColor!=0)
////            outputColor = fairyColor;
////        else if (bulletColor!=0)
////            outputColor = bulletColor;
////        else
////            outputColor = 5'b0; // set this to background later?
////
////        palette_out = outputColor;
//			palette_out = playerColor;
//    end
//
//endmodule
